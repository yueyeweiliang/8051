module INST_EXT(INT_REQ, MONITOR_REQUEST, BREAK_FLAG, INSTR_EXTN, INT_LEVEL, REAL_TIME_ON);
input INT_REQ, MONITOR_REQUEST, BREAK_FLAG;
input  [1:0] INT_LEVEL;
output [2:0] INSTR_EXTN;
input		 REAL_TIME_ON;

reg [2:0] INSTR_EXTN;


always @(INT_REQ or MONITOR_REQUEST or BREAK_FLAG or INT_LEVEL or REAL_TIME_ON) begin
	if (MONITOR_REQUEST ) INSTR_EXTN = 3'b100;
	else if (INT_REQ & ~(BREAK_FLAG & ~REAL_TIME_ON)) 	 INSTR_EXTN = 3'b010;
	else if (BREAK_FLAG & ~|INT_LEVEL) INSTR_EXTN = 3'b001;
	else 				 INSTR_EXTN = 3'b000;
end	


endmodule
